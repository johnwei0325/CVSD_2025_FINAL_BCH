// LUT
// (63, 51) BCH
module GF_06 (
	input [5:0] power,
	output reg [5:0] poly
);
	always @* begin
		case(power)
			6'd-1: poly = 6'd0;
			6'd0: poly = 6'd1;
			6'd1: poly = 6'd2;
			6'd2: poly = 6'd4;
			6'd3: poly = 6'd8;
			6'd4: poly = 6'd16;
			6'd5: poly = 6'd32;
			6'd6: poly = 6'd3;
			6'd7: poly = 6'd6;
			6'd8: poly = 6'd12;
			6'd9: poly = 6'd24;
			6'd10: poly = 6'd48;
			6'd11: poly = 6'd35;
			6'd12: poly = 6'd5;
			6'd13: poly = 6'd10;
			6'd14: poly = 6'd20;
			6'd15: poly = 6'd40;
			6'd16: poly = 6'd19;
			6'd17: poly = 6'd38;
			6'd18: poly = 6'd15;
			6'd19: poly = 6'd30;
			6'd20: poly = 6'd60;
			6'd21: poly = 6'd59;
			6'd22: poly = 6'd53;
			6'd23: poly = 6'd41;
			6'd24: poly = 6'd17;
			6'd25: poly = 6'd34;
			6'd26: poly = 6'd7;
			6'd27: poly = 6'd14;
			6'd28: poly = 6'd28;
			6'd29: poly = 6'd56;
			6'd30: poly = 6'd51;
			6'd31: poly = 6'd37;
			6'd32: poly = 6'd9;
			6'd33: poly = 6'd18;
			6'd34: poly = 6'd36;
			6'd35: poly = 6'd11;
			6'd36: poly = 6'd22;
			6'd37: poly = 6'd44;
			6'd38: poly = 6'd27;
			6'd39: poly = 6'd54;
			6'd40: poly = 6'd47;
			6'd41: poly = 6'd29;
			6'd42: poly = 6'd58;
			6'd43: poly = 6'd55;
			6'd44: poly = 6'd45;
			6'd45: poly = 6'd25;
			6'd46: poly = 6'd50;
			6'd47: poly = 6'd39;
			6'd48: poly = 6'd13;
			6'd49: poly = 6'd26;
			6'd50: poly = 6'd52;
			6'd51: poly = 6'd43;
			6'd52: poly = 6'd21;
			6'd53: poly = 6'd42;
			6'd54: poly = 6'd23;
			6'd55: poly = 6'd46;
			6'd56: poly = 6'd31;
			6'd57: poly = 6'd62;
			6'd58: poly = 6'd63;
			6'd59: poly = 6'd61;
			6'd60: poly = 6'd57;
			6'd61: poly = 6'd49;
			6'd62: poly = 6'd33;
			default: poly = 6'0;
		endcase
	end
endmodule

module GF_06_inv (
	input [5:0] poly,
	output reg [5:0] power
);
	always @* begin
		case(poly)
			6'd0: power = 6'd-1;
			6'd1: power = 6'd0;
			6'd2: power = 6'd1;
			6'd4: power = 6'd2;
			6'd8: power = 6'd3;
			6'd16: power = 6'd4;
			6'd32: power = 6'd5;
			6'd3: power = 6'd6;
			6'd6: power = 6'd7;
			6'd12: power = 6'd8;
			6'd24: power = 6'd9;
			6'd48: power = 6'd10;
			6'd35: power = 6'd11;
			6'd5: power = 6'd12;
			6'd10: power = 6'd13;
			6'd20: power = 6'd14;
			6'd40: power = 6'd15;
			6'd19: power = 6'd16;
			6'd38: power = 6'd17;
			6'd15: power = 6'd18;
			6'd30: power = 6'd19;
			6'd60: power = 6'd20;
			6'd59: power = 6'd21;
			6'd53: power = 6'd22;
			6'd41: power = 6'd23;
			6'd17: power = 6'd24;
			6'd34: power = 6'd25;
			6'd7: power = 6'd26;
			6'd14: power = 6'd27;
			6'd28: power = 6'd28;
			6'd56: power = 6'd29;
			6'd51: power = 6'd30;
			6'd37: power = 6'd31;
			6'd9: power = 6'd32;
			6'd18: power = 6'd33;
			6'd36: power = 6'd34;
			6'd11: power = 6'd35;
			6'd22: power = 6'd36;
			6'd44: power = 6'd37;
			6'd27: power = 6'd38;
			6'd54: power = 6'd39;
			6'd47: power = 6'd40;
			6'd29: power = 6'd41;
			6'd58: power = 6'd42;
			6'd55: power = 6'd43;
			6'd45: power = 6'd44;
			6'd25: power = 6'd45;
			6'd50: power = 6'd46;
			6'd39: power = 6'd47;
			6'd13: power = 6'd48;
			6'd26: power = 6'd49;
			6'd52: power = 6'd50;
			6'd43: power = 6'd51;
			6'd21: power = 6'd52;
			6'd42: power = 6'd53;
			6'd23: power = 6'd54;
			6'd46: power = 6'd55;
			6'd31: power = 6'd56;
			6'd62: power = 6'd57;
			6'd63: power = 6'd58;
			6'd61: power = 6'd59;
			6'd57: power = 6'd60;
			6'd49: power = 6'd61;
			6'd33: power = 6'd62;
            default : power = 6'd63;
		endcase
	end
endmodule

// (255, 239) BCH
module GF_08 (
	input [7:0] power,
	output reg [7:0] poly
);
	always @* begin
        case(power)
            8'd-1: poly = 8'd0;
            8'd0: poly = 8'd1;
            8'd1: poly = 8'd2;
            8'd2: poly = 8'd4;
            8'd3: poly = 8'd8;
            8'd4: poly = 8'd16;
            8'd5: poly = 8'd32;
            8'd6: poly = 8'd64;
            8'd7: poly = 8'd128;
            8'd8: poly = 8'd29;
            8'd9: poly = 8'd58;
            8'd10: poly = 8'd116;
            8'd11: poly = 8'd232;
            8'd12: poly = 8'd205;
            8'd13: poly = 8'd135;
            8'd14: poly = 8'd19;
            8'd15: poly = 8'd38;
            8'd16: poly = 8'd76;
            8'd17: poly = 8'd152;
            8'd18: poly = 8'd45;
            8'd19: poly = 8'd90;
            8'd20: poly = 8'd180;
            8'd21: poly = 8'd117;
            8'd22: poly = 8'd234;
            8'd23: poly = 8'd201;
            8'd24: poly = 8'd143;
            8'd25: poly = 8'd3;
            8'd26: poly = 8'd6;
            8'd27: poly = 8'd12;
            8'd28: poly = 8'd24;
            8'd29: poly = 8'd48;
            8'd30: poly = 8'd96;
            8'd31: poly = 8'd192;
            8'd32: poly = 8'd157;
            8'd33: poly = 8'd39;
            8'd34: poly = 8'd78;
            8'd35: poly = 8'd156;
            8'd36: poly = 8'd37;
            8'd37: poly = 8'd74;
            8'd38: poly = 8'd148;
            8'd39: poly = 8'd53;
            8'd40: poly = 8'd106;
            8'd41: poly = 8'd212;
            8'd42: poly = 8'd181;
            8'd43: poly = 8'd119;
            8'd44: poly = 8'd238;
            8'd45: poly = 8'd193;
            8'd46: poly = 8'd159;
            8'd47: poly = 8'd35;
            8'd48: poly = 8'd70;
            8'd49: poly = 8'd140;
            8'd50: poly = 8'd5;
            8'd51: poly = 8'd10;
            8'd52: poly = 8'd20;
            8'd53: poly = 8'd40;
            8'd54: poly = 8'd80;
            8'd55: poly = 8'd160;
            8'd56: poly = 8'd93;
            8'd57: poly = 8'd186;
            8'd58: poly = 8'd105;
            8'd59: poly = 8'd210;
            8'd60: poly = 8'd185;
            8'd61: poly = 8'd111;
            8'd62: poly = 8'd222;
            8'd63: poly = 8'd161;
            8'd64: poly = 8'd95;
            8'd65: poly = 8'd190;
            8'd66: poly = 8'd97;
            8'd67: poly = 8'd194;
            8'd68: poly = 8'd153;
            8'd69: poly = 8'd47;
            8'd70: poly = 8'd94;
            8'd71: poly = 8'd188;
            8'd72: poly = 8'd101;
            8'd73: poly = 8'd202;
            8'd74: poly = 8'd137;
            8'd75: poly = 8'd15;
            8'd76: poly = 8'd30;
            8'd77: poly = 8'd60;
            8'd78: poly = 8'd120;
            8'd79: poly = 8'd240;
            8'd80: poly = 8'd253;
            8'd81: poly = 8'd231;
            8'd82: poly = 8'd211;
            8'd83: poly = 8'd187;
            8'd84: poly = 8'd107;
            8'd85: poly = 8'd214;
            8'd86: poly = 8'd177;
            8'd87: poly = 8'd127;
            8'd88: poly = 8'd254;
            8'd89: poly = 8'd225;
            8'd90: poly = 8'd223;
            8'd91: poly = 8'd163;
            8'd92: poly = 8'd91;
            8'd93: poly = 8'd182;
            8'd94: poly = 8'd113;
            8'd95: poly = 8'd226;
            8'd96: poly = 8'd217;
            8'd97: poly = 8'd175;
            8'd98: poly = 8'd67;
            8'd99: poly = 8'd134;
            8'd100: poly = 8'd17;
            8'd101: poly = 8'd34;
            8'd102: poly = 8'd68;
            8'd103: poly = 8'd136;
            8'd104: poly = 8'd13;
            8'd105: poly = 8'd26;
            8'd106: poly = 8'd52;
            8'd107: poly = 8'd104;
            8'd108: poly = 8'd208;
            8'd109: poly = 8'd189;
            8'd110: poly = 8'd103;
            8'd111: poly = 8'd206;
            8'd112: poly = 8'd129;
            8'd113: poly = 8'd31;
            8'd114: poly = 8'd62;
            8'd115: poly = 8'd124;
            8'd116: poly = 8'd248;
            8'd117: poly = 8'd237;
            8'd118: poly = 8'd199;
            8'd119: poly = 8'd147;
            8'd120: poly = 8'd59;
            8'd121: poly = 8'd118;
            8'd122: poly = 8'd236;
            8'd123: poly = 8'd197;
            8'd124: poly = 8'd151;
            8'd125: poly = 8'd51;
            8'd126: poly = 8'd102;
            8'd127: poly = 8'd204;
            8'd128: poly = 8'd133;
            8'd129: poly = 8'd23;
            8'd130: poly = 8'd46;
            8'd131: poly = 8'd92;
            8'd132: poly = 8'd184;
            8'd133: poly = 8'd109;
            8'd134: poly = 8'd218;
            8'd135: poly = 8'd169;
            8'd136: poly = 8'd79;
            8'd137: poly = 8'd158;
            8'd138: poly = 8'd33;
            8'd139: poly = 8'd66;
            8'd140: poly = 8'd132;
            8'd141: poly = 8'd21;
            8'd142: poly = 8'd42;
            8'd143: poly = 8'd84;
            8'd144: poly = 8'd168;
            8'd145: poly = 8'd77;
            8'd146: poly = 8'd154;
            8'd147: poly = 8'd41;
            8'd148: poly = 8'd82;
            8'd149: poly = 8'd164;
            8'd150: poly = 8'd85;
            8'd151: poly = 8'd170;
            8'd152: poly = 8'd73;
            8'd153: poly = 8'd146;
            8'd154: poly = 8'd57;
            8'd155: poly = 8'd114;
            8'd156: poly = 8'd228;
            8'd157: poly = 8'd213;
            8'd158: poly = 8'd183;
            8'd159: poly = 8'd115;
            8'd160: poly = 8'd230;
            8'd161: poly = 8'd209;
            8'd162: poly = 8'd191;
            8'd163: poly = 8'd99;
            8'd164: poly = 8'd198;
            8'd165: poly = 8'd145;
            8'd166: poly = 8'd63;
            8'd167: poly = 8'd126;
            8'd168: poly = 8'd252;
            8'd169: poly = 8'd229;
            8'd170: poly = 8'd215;
            8'd171: poly = 8'd179;
            8'd172: poly = 8'd123;
            8'd173: poly = 8'd246;
            8'd174: poly = 8'd241;
            8'd175: poly = 8'd255;
            8'd176: poly = 8'd227;
            8'd177: poly = 8'd219;
            8'd178: poly = 8'd171;
            8'd179: poly = 8'd75;
            8'd180: poly = 8'd150;
            8'd181: poly = 8'd49;
            8'd182: poly = 8'd98;
            8'd183: poly = 8'd196;
            8'd184: poly = 8'd149;
            8'd185: poly = 8'd55;
            8'd186: poly = 8'd110;
            8'd187: poly = 8'd220;
            8'd188: poly = 8'd165;
            8'd189: poly = 8'd87;
            8'd190: poly = 8'd174;
            8'd191: poly = 8'd65;
            8'd192: poly = 8'd130;
            8'd193: poly = 8'd25;
            8'd194: poly = 8'd50;
            8'd195: poly = 8'd100;
            8'd196: poly = 8'd200;
            8'd197: poly = 8'd141;
            8'd198: poly = 8'd7;
            8'd199: poly = 8'd14;
            8'd200: poly = 8'd28;
            8'd201: poly = 8'd56;
            8'd202: poly = 8'd112;
            8'd203: poly = 8'd224;
            8'd204: poly = 8'd221;
            8'd205: poly = 8'd167;
            8'd206: poly = 8'd83;
            8'd207: poly = 8'd166;
            8'd208: poly = 8'd81;
            8'd209: poly = 8'd162;
            8'd210: poly = 8'd89;
            8'd211: poly = 8'd178;
            8'd212: poly = 8'd121;
            8'd213: poly = 8'd242;
            8'd214: poly = 8'd249;
            8'd215: poly = 8'd239;
            8'd216: poly = 8'd195;
            8'd217: poly = 8'd155;
            8'd218: poly = 8'd43;
            8'd219: poly = 8'd86;
            8'd220: poly = 8'd172;
            8'd221: poly = 8'd69;
            8'd222: poly = 8'd138;
            8'd223: poly = 8'd9;
            8'd224: poly = 8'd18;
            8'd225: poly = 8'd36;
            8'd226: poly = 8'd72;
            8'd227: poly = 8'd144;
            8'd228: poly = 8'd61;
            8'd229: poly = 8'd122;
            8'd230: poly = 8'd244;
            8'd231: poly = 8'd245;
            8'd232: poly = 8'd247;
            8'd233: poly = 8'd243;
            8'd234: poly = 8'd251;
            8'd235: poly = 8'd235;
            8'd236: poly = 8'd203;
            8'd237: poly = 8'd139;
            8'd238: poly = 8'd11;
            8'd239: poly = 8'd22;
            8'd240: poly = 8'd44;
            8'd241: poly = 8'd88;
            8'd242: poly = 8'd176;
            8'd243: poly = 8'd125;
            8'd244: poly = 8'd250;
            8'd245: poly = 8'd233;
            8'd246: poly = 8'd207;
            8'd247: poly = 8'd131;
            8'd248: poly = 8'd27;
            8'd249: poly = 8'd54;
            8'd250: poly = 8'd108;
            8'd251: poly = 8'd216;
            8'd252: poly = 8'd173;
            8'd253: poly = 8'd71;
            8'd254: poly = 8'd142;
            default: poly = 8'd0;
        endcase
    end

endmodule

module GF_08_inv (
	input [7:0] poly,
	output reg [7:0] power
);
    always @* begin
        case(poly)
            8'd0: power = 8'd-1;
            8'd1: power = 8'd0;
            8'd2: power = 8'd1;
            8'd4: power = 8'd2;
            8'd8: power = 8'd3;
            8'd16: power = 8'd4;
            8'd32: power = 8'd5;
            8'd64: power = 8'd6;
            8'd128: power = 8'd7;
            8'd29: power = 8'd8;
            8'd58: power = 8'd9;
            8'd116: power = 8'd10;
            8'd232: power = 8'd11;
            8'd205: power = 8'd12;
            8'd135: power = 8'd13;
            8'd19: power = 8'd14;
            8'd38: power = 8'd15;
            8'd76: power = 8'd16;
            8'd152: power = 8'd17;
            8'd45: power = 8'd18;
            8'd90: power = 8'd19;
            8'd180: power = 8'd20;
            8'd117: power = 8'd21;
            8'd234: power = 8'd22;
            8'd201: power = 8'd23;
            8'd143: power = 8'd24;
            8'd3: power = 8'd25;
            8'd6: power = 8'd26;
            8'd12: power = 8'd27;
            8'd24: power = 8'd28;
            8'd48: power = 8'd29;
            8'd96: power = 8'd30;
            8'd192: power = 8'd31;
            8'd157: power = 8'd32;
            8'd39: power = 8'd33;
            8'd78: power = 8'd34;
            8'd156: power = 8'd35;
            8'd37: power = 8'd36;
            8'd74: power = 8'd37;
            8'd148: power = 8'd38;
            8'd53: power = 8'd39;
            8'd106: power = 8'd40;
            8'd212: power = 8'd41;
            8'd181: power = 8'd42;
            8'd119: power = 8'd43;
            8'd238: power = 8'd44;
            8'd193: power = 8'd45;
            8'd159: power = 8'd46;
            8'd35: power = 8'd47;
            8'd70: power = 8'd48;
            8'd140: power = 8'd49;
            8'd5: power = 8'd50;
            8'd10: power = 8'd51;
            8'd20: power = 8'd52;
            8'd40: power = 8'd53;
            8'd80: power = 8'd54;
            8'd160: power = 8'd55;
            8'd93: power = 8'd56;
            8'd186: power = 8'd57;
            8'd105: power = 8'd58;
            8'd210: power = 8'd59;
            8'd185: power = 8'd60;
            8'd111: power = 8'd61;
            8'd222: power = 8'd62;
            8'd161: power = 8'd63;
            8'd95: power = 8'd64;
            8'd190: power = 8'd65;
            8'd97: power = 8'd66;
            8'd194: power = 8'd67;
            8'd153: power = 8'd68;
            8'd47: power = 8'd69;
            8'd94: power = 8'd70;
            8'd188: power = 8'd71;
            8'd101: power = 8'd72;
            8'd202: power = 8'd73;
            8'd137: power = 8'd74;
            8'd15: power = 8'd75;
            8'd30: power = 8'd76;
            8'd60: power = 8'd77;
            8'd120: power = 8'd78;
            8'd240: power = 8'd79;
            8'd253: power = 8'd80;
            8'd231: power = 8'd81;
            8'd211: power = 8'd82;
            8'd187: power = 8'd83;
            8'd107: power = 8'd84;
            8'd214: power = 8'd85;
            8'd177: power = 8'd86;
            8'd127: power = 8'd87;
            8'd254: power = 8'd88;
            8'd225: power = 8'd89;
            8'd223: power = 8'd90;
            8'd163: power = 8'd91;
            8'd91: power = 8'd92;
            8'd182: power = 8'd93;
            8'd113: power = 8'd94;
            8'd226: power = 8'd95;
            8'd217: power = 8'd96;
            8'd175: power = 8'd97;
            8'd67: power = 8'd98;
            8'd134: power = 8'd99;
            8'd17: power = 8'd100;
            8'd34: power = 8'd101;
            8'd68: power = 8'd102;
            8'd136: power = 8'd103;
            8'd13: power = 8'd104;
            8'd26: power = 8'd105;
            8'd52: power = 8'd106;
            8'd104: power = 8'd107;
            8'd208: power = 8'd108;
            8'd189: power = 8'd109;
            8'd103: power = 8'd110;
            8'd206: power = 8'd111;
            8'd129: power = 8'd112;
            8'd31: power = 8'd113;
            8'd62: power = 8'd114;
            8'd124: power = 8'd115;
            8'd248: power = 8'd116;
            8'd237: power = 8'd117;
            8'd199: power = 8'd118;
            8'd147: power = 8'd119;
            8'd59: power = 8'd120;
            8'd118: power = 8'd121;
            8'd236: power = 8'd122;
            8'd197: power = 8'd123;
            8'd151: power = 8'd124;
            8'd51: power = 8'd125;
            8'd102: power = 8'd126;
            8'd204: power = 8'd127;
            8'd133: power = 8'd128;
            8'd23: power = 8'd129;
            8'd46: power = 8'd130;
            8'd92: power = 8'd131;
            8'd184: power = 8'd132;
            8'd109: power = 8'd133;
            8'd218: power = 8'd134;
            8'd169: power = 8'd135;
            8'd79: power = 8'd136;
            8'd158: power = 8'd137;
            8'd33: power = 8'd138;
            8'd66: power = 8'd139;
            8'd132: power = 8'd140;
            8'd21: power = 8'd141;
            8'd42: power = 8'd142;
            8'd84: power = 8'd143;
            8'd168: power = 8'd144;
            8'd77: power = 8'd145;
            8'd154: power = 8'd146;
            8'd41: power = 8'd147;
            8'd82: power = 8'd148;
            8'd164: power = 8'd149;
            8'd85: power = 8'd150;
            8'd170: power = 8'd151;
            8'd73: power = 8'd152;
            8'd146: power = 8'd153;
            8'd57: power = 8'd154;
            8'd114: power = 8'd155;
            8'd228: power = 8'd156;
            8'd213: power = 8'd157;
            8'd183: power = 8'd158;
            8'd115: power = 8'd159;
            8'd230: power = 8'd160;
            8'd209: power = 8'd161;
            8'd191: power = 8'd162;
            8'd99: power = 8'd163;
            8'd198: power = 8'd164;
            8'd145: power = 8'd165;
            8'd63: power = 8'd166;
            8'd126: power = 8'd167;
            8'd252: power = 8'd168;
            8'd229: power = 8'd169;
            8'd215: power = 8'd170;
            8'd179: power = 8'd171;
            8'd123: power = 8'd172;
            8'd246: power = 8'd173;
            8'd241: power = 8'd174;
            8'd255: power = 8'd175;
            8'd227: power = 8'd176;
            8'd219: power = 8'd177;
            8'd171: power = 8'd178;
            8'd75: power = 8'd179;
            8'd150: power = 8'd180;
            8'd49: power = 8'd181;
            8'd98: power = 8'd182;
            8'd196: power = 8'd183;
            8'd149: power = 8'd184;
            8'd55: power = 8'd185;
            8'd110: power = 8'd186;
            8'd220: power = 8'd187;
            8'd165: power = 8'd188;
            8'd87: power = 8'd189;
            8'd174: power = 8'd190;
            8'd65: power = 8'd191;
            8'd130: power = 8'd192;
            8'd25: power = 8'd193;
            8'd50: power = 8'd194;
            8'd100: power = 8'd195;
            8'd200: power = 8'd196;
            8'd141: power = 8'd197;
            8'd7: power = 8'd198;
            8'd14: power = 8'd199;
            8'd28: power = 8'd200;
            8'd56: power = 8'd201;
            8'd112: power = 8'd202;
            8'd224: power = 8'd203;
            8'd221: power = 8'd204;
            8'd167: power = 8'd205;
            8'd83: power = 8'd206;
            8'd166: power = 8'd207;
            8'd81: power = 8'd208;
            8'd162: power = 8'd209;
            8'd89: power = 8'd210;
            8'd178: power = 8'd211;
            8'd121: power = 8'd212;
            8'd242: power = 8'd213;
            8'd249: power = 8'd214;
            8'd239: power = 8'd215;
            8'd195: power = 8'd216;
            8'd155: power = 8'd217;
            8'd43: power = 8'd218;
            8'd86: power = 8'd219;
            8'd172: power = 8'd220;
            8'd69: power = 8'd221;
            8'd138: power = 8'd222;
            8'd9: power = 8'd223;
            8'd18: power = 8'd224;
            8'd36: power = 8'd225;
            8'd72: power = 8'd226;
            8'd144: power = 8'd227;
            8'd61: power = 8'd228;
            8'd122: power = 8'd229;
            8'd244: power = 8'd230;
            8'd245: power = 8'd231;
            8'd247: power = 8'd232;
            8'd243: power = 8'd233;
            8'd251: power = 8'd234;
            8'd235: power = 8'd235;
            8'd203: power = 8'd236;
            8'd139: power = 8'd237;
            8'd11: power = 8'd238;
            8'd22: power = 8'd239;
            8'd44: power = 8'd240;
            8'd88: power = 8'd241;
            8'd176: power = 8'd242;
            8'd125: power = 8'd243;
            8'd250: power = 8'd244;
            8'd233: power = 8'd245;
            8'd207: power = 8'd246;
            8'd131: power = 8'd247;
            8'd27: power = 8'd248;
            8'd54: power = 8'd249;
            8'd108: power = 8'd250;
            8'd216: power = 8'd251;
            8'd173: power = 8'd252;
            8'd71: power = 8'd253;
            8'd142: power = 8'd254;
            default: power = 8'd255;
        endcase
    end
endmodule

// (1023, 983) BCH
module GF_10 (
	input [9:0] power,
	output reg [9:0] poly
);
	always @* begin
        case(power)
            10'd-1: poly = 10'd0;
            10'd0: poly = 10'd1;
            10'd1: poly = 10'd2;
            10'd2: poly = 10'd4;
            10'd3: poly = 10'd8;
            10'd4: poly = 10'd16;
            10'd5: poly = 10'd32;
            10'd6: poly = 10'd64;
            10'd7: poly = 10'd128;
            10'd8: poly = 10'd256;
            10'd9: poly = 10'd512;
            10'd10: poly = 10'd9;
            10'd11: poly = 10'd18;
            10'd12: poly = 10'd36;
            10'd13: poly = 10'd72;
            10'd14: poly = 10'd144;
            10'd15: poly = 10'd288;
            10'd16: poly = 10'd576;
            10'd17: poly = 10'd137;
            10'd18: poly = 10'd274;
            10'd19: poly = 10'd548;
            10'd20: poly = 10'd65;
            10'd21: poly = 10'd130;
            10'd22: poly = 10'd260;
            10'd23: poly = 10'd520;
            10'd24: poly = 10'd25;
            10'd25: poly = 10'd50;
            10'd26: poly = 10'd100;
            10'd27: poly = 10'd200;
            10'd28: poly = 10'd400;
            10'd29: poly = 10'd800;
            10'd30: poly = 10'd585;
            10'd31: poly = 10'd155;
            10'd32: poly = 10'd310;
            10'd33: poly = 10'd620;
            10'd34: poly = 10'd209;
            10'd35: poly = 10'd418;
            10'd36: poly = 10'd836;
            10'd37: poly = 10'd641;
            10'd38: poly = 10'd267;
            10'd39: poly = 10'd534;
            10'd40: poly = 10'd37;
            10'd41: poly = 10'd74;
            10'd42: poly = 10'd148;
            10'd43: poly = 10'd296;
            10'd44: poly = 10'd592;
            10'd45: poly = 10'd169;
            10'd46: poly = 10'd338;
            10'd47: poly = 10'd676;
            10'd48: poly = 10'd321;
            10'd49: poly = 10'd642;
            10'd50: poly = 10'd269;
            10'd51: poly = 10'd538;
            10'd52: poly = 10'd61;
            10'd53: poly = 10'd122;
            10'd54: poly = 10'd244;
            10'd55: poly = 10'd488;
            10'd56: poly = 10'd976;
            10'd57: poly = 10'd937;
            10'd58: poly = 10'd859;
            10'd59: poly = 10'd703;
            10'd60: poly = 10'd375;
            10'd61: poly = 10'd750;
            10'd62: poly = 10'd469;
            10'd63: poly = 10'd938;
            10'd64: poly = 10'd861;
            10'd65: poly = 10'd691;
            10'd66: poly = 10'd367;
            10'd67: poly = 10'd734;
            10'd68: poly = 10'd437;
            10'd69: poly = 10'd874;
            10'd70: poly = 10'd733;
            10'd71: poly = 10'd435;
            10'd72: poly = 10'd870;
            10'd73: poly = 10'd709;
            10'd74: poly = 10'd387;
            10'd75: poly = 10'd774;
            10'd76: poly = 10'd517;
            10'd77: poly = 10'd3;
            10'd78: poly = 10'd6;
            10'd79: poly = 10'd12;
            10'd80: poly = 10'd24;
            10'd81: poly = 10'd48;
            10'd82: poly = 10'd96;
            10'd83: poly = 10'd192;
            10'd84: poly = 10'd384;
            10'd85: poly = 10'd768;
            10'd86: poly = 10'd521;
            10'd87: poly = 10'd27;
            10'd88: poly = 10'd54;
            10'd89: poly = 10'd108;
            10'd90: poly = 10'd216;
            10'd91: poly = 10'd432;
            10'd92: poly = 10'd864;
            10'd93: poly = 10'd713;
            10'd94: poly = 10'd411;
            10'd95: poly = 10'd822;
            10'd96: poly = 10'd613;
            10'd97: poly = 10'd195;
            10'd98: poly = 10'd390;
            10'd99: poly = 10'd780;
            10'd100: poly = 10'd529;
            10'd101: poly = 10'd43;
            10'd102: poly = 10'd86;
            10'd103: poly = 10'd172;
            10'd104: poly = 10'd344;
            10'd105: poly = 10'd688;
            10'd106: poly = 10'd361;
            10'd107: poly = 10'd722;
            10'd108: poly = 10'd429;
            10'd109: poly = 10'd858;
            10'd110: poly = 10'd701;
            10'd111: poly = 10'd371;
            10'd112: poly = 10'd742;
            10'd113: poly = 10'd453;
            10'd114: poly = 10'd906;
            10'd115: poly = 10'd797;
            10'd116: poly = 10'd563;
            10'd117: poly = 10'd111;
            10'd118: poly = 10'd222;
            10'd119: poly = 10'd444;
            10'd120: poly = 10'd888;
            10'd121: poly = 10'd761;
            10'd122: poly = 10'd507;
            10'd123: poly = 10'd1014;
            10'd124: poly = 10'd997;
            10'd125: poly = 10'd963;
            10'd126: poly = 10'd911;
            10'd127: poly = 10'd791;
            10'd128: poly = 10'd551;
            10'd129: poly = 10'd71;
            10'd130: poly = 10'd142;
            10'd131: poly = 10'd284;
            10'd132: poly = 10'd568;
            10'd133: poly = 10'd121;
            10'd134: poly = 10'd242;
            10'd135: poly = 10'd484;
            10'd136: poly = 10'd968;
            10'd137: poly = 10'd921;
            10'd138: poly = 10'd827;
            10'd139: poly = 10'd639;
            10'd140: poly = 10'd247;
            10'd141: poly = 10'd494;
            10'd142: poly = 10'd988;
            10'd143: poly = 10'd945;
            10'd144: poly = 10'd875;
            10'd145: poly = 10'd735;
            10'd146: poly = 10'd439;
            10'd147: poly = 10'd878;
            10'd148: poly = 10'd725;
            10'd149: poly = 10'd419;
            10'd150: poly = 10'd838;
            10'd151: poly = 10'd645;
            10'd152: poly = 10'd259;
            10'd153: poly = 10'd518;
            10'd154: poly = 10'd5;
            10'd155: poly = 10'd10;
            10'd156: poly = 10'd20;
            10'd157: poly = 10'd40;
            10'd158: poly = 10'd80;
            10'd159: poly = 10'd160;
            10'd160: poly = 10'd320;
            10'd161: poly = 10'd640;
            10'd162: poly = 10'd265;
            10'd163: poly = 10'd530;
            10'd164: poly = 10'd45;
            10'd165: poly = 10'd90;
            10'd166: poly = 10'd180;
            10'd167: poly = 10'd360;
            10'd168: poly = 10'd720;
            10'd169: poly = 10'd425;
            10'd170: poly = 10'd850;
            10'd171: poly = 10'd685;
            10'd172: poly = 10'd339;
            10'd173: poly = 10'd678;
            10'd174: poly = 10'd325;
            10'd175: poly = 10'd650;
            10'd176: poly = 10'd285;
            10'd177: poly = 10'd570;
            10'd178: poly = 10'd125;
            10'd179: poly = 10'd250;
            10'd180: poly = 10'd500;
            10'd181: poly = 10'd1000;
            10'd182: poly = 10'd985;
            10'd183: poly = 10'd955;
            10'd184: poly = 10'd895;
            10'd185: poly = 10'd759;
            10'd186: poly = 10'd487;
            10'd187: poly = 10'd974;
            10'd188: poly = 10'd917;
            10'd189: poly = 10'd803;
            10'd190: poly = 10'd591;
            10'd191: poly = 10'd151;
            10'd192: poly = 10'd302;
            10'd193: poly = 10'd604;
            10'd194: poly = 10'd177;
            10'd195: poly = 10'd354;
            10'd196: poly = 10'd708;
            10'd197: poly = 10'd385;
            10'd198: poly = 10'd770;
            10'd199: poly = 10'd525;
            10'd200: poly = 10'd19;
            10'd201: poly = 10'd38;
            10'd202: poly = 10'd76;
            10'd203: poly = 10'd152;
            10'd204: poly = 10'd304;
            10'd205: poly = 10'd608;
            10'd206: poly = 10'd201;
            10'd207: poly = 10'd402;
            10'd208: poly = 10'd804;
            10'd209: poly = 10'd577;
            10'd210: poly = 10'd139;
            10'd211: poly = 10'd278;
            10'd212: poly = 10'd556;
            10'd213: poly = 10'd81;
            10'd214: poly = 10'd162;
            10'd215: poly = 10'd324;
            10'd216: poly = 10'd648;
            10'd217: poly = 10'd281;
            10'd218: poly = 10'd562;
            10'd219: poly = 10'd109;
            10'd220: poly = 10'd218;
            10'd221: poly = 10'd436;
            10'd222: poly = 10'd872;
            10'd223: poly = 10'd729;
            10'd224: poly = 10'd443;
            10'd225: poly = 10'd886;
            10'd226: poly = 10'd741;
            10'd227: poly = 10'd451;
            10'd228: poly = 10'd902;
            10'd229: poly = 10'd773;
            10'd230: poly = 10'd515;
            10'd231: poly = 10'd15;
            10'd232: poly = 10'd30;
            10'd233: poly = 10'd60;
            10'd234: poly = 10'd120;
            10'd235: poly = 10'd240;
            10'd236: poly = 10'd480;
            10'd237: poly = 10'd960;
            10'd238: poly = 10'd905;
            10'd239: poly = 10'd795;
            10'd240: poly = 10'd575;
            10'd241: poly = 10'd119;
            10'd242: poly = 10'd238;
            10'd243: poly = 10'd476;
            10'd244: poly = 10'd952;
            10'd245: poly = 10'd889;
            10'd246: poly = 10'd763;
            10'd247: poly = 10'd511;
            10'd248: poly = 10'd1022;
            10'd249: poly = 10'd1013;
            10'd250: poly = 10'd995;
            10'd251: poly = 10'd975;
            10'd252: poly = 10'd919;
            10'd253: poly = 10'd807;
            10'd254: poly = 10'd583;
            10'd255: poly = 10'd135;
            10'd256: poly = 10'd270;
            10'd257: poly = 10'd540;
            10'd258: poly = 10'd49;
            10'd259: poly = 10'd98;
            10'd260: poly = 10'd196;
            10'd261: poly = 10'd392;
            10'd262: poly = 10'd784;
            10'd263: poly = 10'd553;
            10'd264: poly = 10'd91;
            10'd265: poly = 10'd182;
            10'd266: poly = 10'd364;
            10'd267: poly = 10'd728;
            10'd268: poly = 10'd441;
            10'd269: poly = 10'd882;
            10'd270: poly = 10'd749;
            10'd271: poly = 10'd467;
            10'd272: poly = 10'd934;
            10'd273: poly = 10'd837;
            10'd274: poly = 10'd643;
            10'd275: poly = 10'd271;
            10'd276: poly = 10'd542;
            10'd277: poly = 10'd53;
            10'd278: poly = 10'd106;
            10'd279: poly = 10'd212;
            10'd280: poly = 10'd424;
            10'd281: poly = 10'd848;
            10'd282: poly = 10'd681;
            10'd283: poly = 10'd347;
            10'd284: poly = 10'd694;
            10'd285: poly = 10'd357;
            10'd286: poly = 10'd714;
            10'd287: poly = 10'd413;
            10'd288: poly = 10'd826;
            10'd289: poly = 10'd637;
            10'd290: poly = 10'd243;
            10'd291: poly = 10'd486;
            10'd292: poly = 10'd972;
            10'd293: poly = 10'd913;
            10'd294: poly = 10'd811;
            10'd295: poly = 10'd607;
            10'd296: poly = 10'd183;
            10'd297: poly = 10'd366;
            10'd298: poly = 10'd732;
            10'd299: poly = 10'd433;
            10'd300: poly = 10'd866;
            10'd301: poly = 10'd717;
            10'd302: poly = 10'd403;
            10'd303: poly = 10'd806;
            10'd304: poly = 10'd581;
            10'd305: poly = 10'd131;
            10'd306: poly = 10'd262;
            10'd307: poly = 10'd524;
            10'd308: poly = 10'd17;
            10'd309: poly = 10'd34;
            10'd310: poly = 10'd68;
            10'd311: poly = 10'd136;
            10'd312: poly = 10'd272;
            10'd313: poly = 10'd544;
            10'd314: poly = 10'd73;
            10'd315: poly = 10'd146;
            10'd316: poly = 10'd292;
            10'd317: poly = 10'd584;
            10'd318: poly = 10'd153;
            10'd319: poly = 10'd306;
            10'd320: poly = 10'd612;
            10'd321: poly = 10'd193;
            10'd322: poly = 10'd386;
            10'd323: poly = 10'd772;
            10'd324: poly = 10'd513;
            10'd325: poly = 10'd11;
            10'd326: poly = 10'd22;
            10'd327: poly = 10'd44;
            10'd328: poly = 10'd88;
            10'd329: poly = 10'd176;
            10'd330: poly = 10'd352;
            10'd331: poly = 10'd704;
            10'd332: poly = 10'd393;
            10'd333: poly = 10'd786;
            10'd334: poly = 10'd557;
            10'd335: poly = 10'd83;
            10'd336: poly = 10'd166;
            10'd337: poly = 10'd332;
            10'd338: poly = 10'd664;
            10'd339: poly = 10'd313;
            10'd340: poly = 10'd626;
            10'd341: poly = 10'd237;
            10'd342: poly = 10'd474;
            10'd343: poly = 10'd948;
            10'd344: poly = 10'd865;
            10'd345: poly = 10'd715;
            10'd346: poly = 10'd415;
            10'd347: poly = 10'd830;
            10'd348: poly = 10'd629;
            10'd349: poly = 10'd227;
            10'd350: poly = 10'd454;
            10'd351: poly = 10'd908;
            10'd352: poly = 10'd785;
            10'd353: poly = 10'd555;
            10'd354: poly = 10'd95;
            10'd355: poly = 10'd190;
            10'd356: poly = 10'd380;
            10'd357: poly = 10'd760;
            10'd358: poly = 10'd505;
            10'd359: poly = 10'd1010;
            10'd360: poly = 10'd1005;
            10'd361: poly = 10'd979;
            10'd362: poly = 10'd943;
            10'd363: poly = 10'd855;
            10'd364: poly = 10'd679;
            10'd365: poly = 10'd327;
            10'd366: poly = 10'd654;
            10'd367: poly = 10'd277;
            10'd368: poly = 10'd554;
            10'd369: poly = 10'd93;
            10'd370: poly = 10'd186;
            10'd371: poly = 10'd372;
            10'd372: poly = 10'd744;
            10'd373: poly = 10'd473;
            10'd374: poly = 10'd946;
            10'd375: poly = 10'd877;
            10'd376: poly = 10'd723;
            10'd377: poly = 10'd431;
            10'd378: poly = 10'd862;
            10'd379: poly = 10'd693;
            10'd380: poly = 10'd355;
            10'd381: poly = 10'd710;
            10'd382: poly = 10'd389;
            10'd383: poly = 10'd778;
            10'd384: poly = 10'd541;
            10'd385: poly = 10'd51;
            10'd386: poly = 10'd102;
            10'd387: poly = 10'd204;
            10'd388: poly = 10'd408;
            10'd389: poly = 10'd816;
            10'd390: poly = 10'd617;
            10'd391: poly = 10'd219;
            10'd392: poly = 10'd438;
            10'd393: poly = 10'd876;
            10'd394: poly = 10'd721;
            10'd395: poly = 10'd427;
            10'd396: poly = 10'd854;
            10'd397: poly = 10'd677;
            10'd398: poly = 10'd323;
            10'd399: poly = 10'd646;
            10'd400: poly = 10'd261;
            10'd401: poly = 10'd522;
            10'd402: poly = 10'd29;
            10'd403: poly = 10'd58;
            10'd404: poly = 10'd116;
            10'd405: poly = 10'd232;
            10'd406: poly = 10'd464;
            10'd407: poly = 10'd928;
            10'd408: poly = 10'd841;
            10'd409: poly = 10'd667;
            10'd410: poly = 10'd319;
            10'd411: poly = 10'd638;
            10'd412: poly = 10'd245;
            10'd413: poly = 10'd490;
            10'd414: poly = 10'd980;
            10'd415: poly = 10'd929;
            10'd416: poly = 10'd843;
            10'd417: poly = 10'd671;
            10'd418: poly = 10'd311;
            10'd419: poly = 10'd622;
            10'd420: poly = 10'd213;
            10'd421: poly = 10'd426;
            10'd422: poly = 10'd852;
            10'd423: poly = 10'd673;
            10'd424: poly = 10'd331;
            10'd425: poly = 10'd662;
            10'd426: poly = 10'd293;
            10'd427: poly = 10'd586;
            10'd428: poly = 10'd157;
            10'd429: poly = 10'd314;
            10'd430: poly = 10'd628;
            10'd431: poly = 10'd225;
            10'd432: poly = 10'd450;
            10'd433: poly = 10'd900;
            10'd434: poly = 10'd769;
            10'd435: poly = 10'd523;
            10'd436: poly = 10'd31;
            10'd437: poly = 10'd62;
            10'd438: poly = 10'd124;
            10'd439: poly = 10'd248;
            10'd440: poly = 10'd496;
            10'd441: poly = 10'd992;
            10'd442: poly = 10'd969;
            10'd443: poly = 10'd923;
            10'd444: poly = 10'd831;
            10'd445: poly = 10'd631;
            10'd446: poly = 10'd231;
            10'd447: poly = 10'd462;
            10'd448: poly = 10'd924;
            10'd449: poly = 10'd817;
            10'd450: poly = 10'd619;
            10'd451: poly = 10'd223;
            10'd452: poly = 10'd446;
            10'd453: poly = 10'd892;
            10'd454: poly = 10'd753;
            10'd455: poly = 10'd491;
            10'd456: poly = 10'd982;
            10'd457: poly = 10'd933;
            10'd458: poly = 10'd835;
            10'd459: poly = 10'd655;
            10'd460: poly = 10'd279;
            10'd461: poly = 10'd558;
            10'd462: poly = 10'd85;
            10'd463: poly = 10'd170;
            10'd464: poly = 10'd340;
            10'd465: poly = 10'd680;
            10'd466: poly = 10'd345;
            10'd467: poly = 10'd690;
            10'd468: poly = 10'd365;
            10'd469: poly = 10'd730;
            10'd470: poly = 10'd445;
            10'd471: poly = 10'd890;
            10'd472: poly = 10'd765;
            10'd473: poly = 10'd499;
            10'd474: poly = 10'd998;
            10'd475: poly = 10'd965;
            10'd476: poly = 10'd899;
            10'd477: poly = 10'd783;
            10'd478: poly = 10'd535;
            10'd479: poly = 10'd39;
            10'd480: poly = 10'd78;
            10'd481: poly = 10'd156;
            10'd482: poly = 10'd312;
            10'd483: poly = 10'd624;
            10'd484: poly = 10'd233;
            10'd485: poly = 10'd466;
            10'd486: poly = 10'd932;
            10'd487: poly = 10'd833;
            10'd488: poly = 10'd651;
            10'd489: poly = 10'd287;
            10'd490: poly = 10'd574;
            10'd491: poly = 10'd117;
            10'd492: poly = 10'd234;
            10'd493: poly = 10'd468;
            10'd494: poly = 10'd936;
            10'd495: poly = 10'd857;
            10'd496: poly = 10'd699;
            10'd497: poly = 10'd383;
            10'd498: poly = 10'd766;
            10'd499: poly = 10'd501;
            10'd500: poly = 10'd1002;
            10'd501: poly = 10'd989;
            10'd502: poly = 10'd947;
            10'd503: poly = 10'd879;
            10'd504: poly = 10'd727;
            10'd505: poly = 10'd423;
            10'd506: poly = 10'd846;
            10'd507: poly = 10'd661;
            10'd508: poly = 10'd291;
            10'd509: poly = 10'd582;
            10'd510: poly = 10'd133;
            10'd511: poly = 10'd266;
            10'd512: poly = 10'd532;
            10'd513: poly = 10'd33;
            10'd514: poly = 10'd66;
            10'd515: poly = 10'd132;
            10'd516: poly = 10'd264;
            10'd517: poly = 10'd528;
            10'd518: poly = 10'd41;
            10'd519: poly = 10'd82;
            10'd520: poly = 10'd164;
            10'd521: poly = 10'd328;
            10'd522: poly = 10'd656;
            10'd523: poly = 10'd297;
            10'd524: poly = 10'd594;
            10'd525: poly = 10'd173;
            10'd526: poly = 10'd346;
            10'd527: poly = 10'd692;
            10'd528: poly = 10'd353;
            10'd529: poly = 10'd706;
            10'd530: poly = 10'd397;
            10'd531: poly = 10'd794;
            10'd532: poly = 10'd573;
            10'd533: poly = 10'd115;
            10'd534: poly = 10'd230;
            10'd535: poly = 10'd460;
            10'd536: poly = 10'd920;
            10'd537: poly = 10'd825;
            10'd538: poly = 10'd635;
            10'd539: poly = 10'd255;
            10'd540: poly = 10'd510;
            10'd541: poly = 10'd1020;
            10'd542: poly = 10'd1009;
            10'd543: poly = 10'd1003;
            10'd544: poly = 10'd991;
            10'd545: poly = 10'd951;
            10'd546: poly = 10'd871;
            10'd547: poly = 10'd711;
            10'd548: poly = 10'd391;
            10'd549: poly = 10'd782;
            10'd550: poly = 10'd533;
            10'd551: poly = 10'd35;
            10'd552: poly = 10'd70;
            10'd553: poly = 10'd140;
            10'd554: poly = 10'd280;
            10'd555: poly = 10'd560;
            10'd556: poly = 10'd105;
            10'd557: poly = 10'd210;
            10'd558: poly = 10'd420;
            10'd559: poly = 10'd840;
            10'd560: poly = 10'd665;
            10'd561: poly = 10'd315;
            10'd562: poly = 10'd630;
            10'd563: poly = 10'd229;
            10'd564: poly = 10'd458;
            10'd565: poly = 10'd916;
            10'd566: poly = 10'd801;
            10'd567: poly = 10'd587;
            10'd568: poly = 10'd159;
            10'd569: poly = 10'd318;
            10'd570: poly = 10'd636;
            10'd571: poly = 10'd241;
            10'd572: poly = 10'd482;
            10'd573: poly = 10'd964;
            10'd574: poly = 10'd897;
            10'd575: poly = 10'd779;
            10'd576: poly = 10'd543;
            10'd577: poly = 10'd55;
            10'd578: poly = 10'd110;
            10'd579: poly = 10'd220;
            10'd580: poly = 10'd440;
            10'd581: poly = 10'd880;
            10'd582: poly = 10'd745;
            10'd583: poly = 10'd475;
            10'd584: poly = 10'd950;
            10'd585: poly = 10'd869;
            10'd586: poly = 10'd707;
            10'd587: poly = 10'd399;
            10'd588: poly = 10'd798;
            10'd589: poly = 10'd565;
            10'd590: poly = 10'd99;
            10'd591: poly = 10'd198;
            10'd592: poly = 10'd396;
            10'd593: poly = 10'd792;
            10'd594: poly = 10'd569;
            10'd595: poly = 10'd123;
            10'd596: poly = 10'd246;
            10'd597: poly = 10'd492;
            10'd598: poly = 10'd984;
            10'd599: poly = 10'd953;
            10'd600: poly = 10'd891;
            10'd601: poly = 10'd767;
            10'd602: poly = 10'd503;
            10'd603: poly = 10'd1006;
            10'd604: poly = 10'd981;
            10'd605: poly = 10'd931;
            10'd606: poly = 10'd847;
            10'd607: poly = 10'd663;
            10'd608: poly = 10'd295;
            10'd609: poly = 10'd590;
            10'd610: poly = 10'd149;
            10'd611: poly = 10'd298;
            10'd612: poly = 10'd596;
            10'd613: poly = 10'd161;
            10'd614: poly = 10'd322;
            10'd615: poly = 10'd644;
            10'd616: poly = 10'd257;
            10'd617: poly = 10'd514;
            10'd618: poly = 10'd13;
            10'd619: poly = 10'd26;
            10'd620: poly = 10'd52;
            10'd621: poly = 10'd104;
            10'd622: poly = 10'd208;
            10'd623: poly = 10'd416;
            10'd624: poly = 10'd832;
            10'd625: poly = 10'd649;
            10'd626: poly = 10'd283;
            10'd627: poly = 10'd566;
            10'd628: poly = 10'd101;
            10'd629: poly = 10'd202;
            10'd630: poly = 10'd404;
            10'd631: poly = 10'd808;
            10'd632: poly = 10'd601;
            10'd633: poly = 10'd187;
            10'd634: poly = 10'd374;
            10'd635: poly = 10'd748;
            10'd636: poly = 10'd465;
            10'd637: poly = 10'd930;
            10'd638: poly = 10'd845;
            10'd639: poly = 10'd659;
            10'd640: poly = 10'd303;
            10'd641: poly = 10'd606;
            10'd642: poly = 10'd181;
            10'd643: poly = 10'd362;
            10'd644: poly = 10'd724;
            10'd645: poly = 10'd417;
            10'd646: poly = 10'd834;
            10'd647: poly = 10'd653;
            10'd648: poly = 10'd275;
            10'd649: poly = 10'd550;
            10'd650: poly = 10'd69;
            10'd651: poly = 10'd138;
            10'd652: poly = 10'd276;
            10'd653: poly = 10'd552;
            10'd654: poly = 10'd89;
            10'd655: poly = 10'd178;
            10'd656: poly = 10'd356;
            10'd657: poly = 10'd712;
            10'd658: poly = 10'd409;
            10'd659: poly = 10'd818;
            10'd660: poly = 10'd621;
            10'd661: poly = 10'd211;
            10'd662: poly = 10'd422;
            10'd663: poly = 10'd844;
            10'd664: poly = 10'd657;
            10'd665: poly = 10'd299;
            10'd666: poly = 10'd598;
            10'd667: poly = 10'd165;
            10'd668: poly = 10'd330;
            10'd669: poly = 10'd660;
            10'd670: poly = 10'd289;
            10'd671: poly = 10'd578;
            10'd672: poly = 10'd141;
            10'd673: poly = 10'd282;
            10'd674: poly = 10'd564;
            10'd675: poly = 10'd97;
            10'd676: poly = 10'd194;
            10'd677: poly = 10'd388;
            10'd678: poly = 10'd776;
            10'd679: poly = 10'd537;
            10'd680: poly = 10'd59;
            10'd681: poly = 10'd118;
            10'd682: poly = 10'd236;
            10'd683: poly = 10'd472;
            10'd684: poly = 10'd944;
            10'd685: poly = 10'd873;
            10'd686: poly = 10'd731;
            10'd687: poly = 10'd447;
            10'd688: poly = 10'd894;
            10'd689: poly = 10'd757;
            10'd690: poly = 10'd483;
            10'd691: poly = 10'd966;
            10'd692: poly = 10'd901;
            10'd693: poly = 10'd771;
            10'd694: poly = 10'd527;
            10'd695: poly = 10'd23;
            10'd696: poly = 10'd46;
            10'd697: poly = 10'd92;
            10'd698: poly = 10'd184;
            10'd699: poly = 10'd368;
            10'd700: poly = 10'd736;
            10'd701: poly = 10'd457;
            10'd702: poly = 10'd914;
            10'd703: poly = 10'd813;
            10'd704: poly = 10'd595;
            10'd705: poly = 10'd175;
            10'd706: poly = 10'd350;
            10'd707: poly = 10'd700;
            10'd708: poly = 10'd369;
            10'd709: poly = 10'd738;
            10'd710: poly = 10'd461;
            10'd711: poly = 10'd922;
            10'd712: poly = 10'd829;
            10'd713: poly = 10'd627;
            10'd714: poly = 10'd239;
            10'd715: poly = 10'd478;
            10'd716: poly = 10'd956;
            10'd717: poly = 10'd881;
            10'd718: poly = 10'd747;
            10'd719: poly = 10'd479;
            10'd720: poly = 10'd958;
            10'd721: poly = 10'd885;
            10'd722: poly = 10'd739;
            10'd723: poly = 10'd463;
            10'd724: poly = 10'd926;
            10'd725: poly = 10'd821;
            10'd726: poly = 10'd611;
            10'd727: poly = 10'd207;
            10'd728: poly = 10'd414;
            10'd729: poly = 10'd828;
            10'd730: poly = 10'd625;
            10'd731: poly = 10'd235;
            10'd732: poly = 10'd470;
            10'd733: poly = 10'd940;
            10'd734: poly = 10'd849;
            10'd735: poly = 10'd683;
            10'd736: poly = 10'd351;
            10'd737: poly = 10'd702;
            10'd738: poly = 10'd373;
            10'd739: poly = 10'd746;
            10'd740: poly = 10'd477;
            10'd741: poly = 10'd954;
            10'd742: poly = 10'd893;
            10'd743: poly = 10'd755;
            10'd744: poly = 10'd495;
            10'd745: poly = 10'd990;
            10'd746: poly = 10'd949;
            10'd747: poly = 10'd867;
            10'd748: poly = 10'd719;
            10'd749: poly = 10'd407;
            10'd750: poly = 10'd814;
            10'd751: poly = 10'd597;
            10'd752: poly = 10'd163;
            10'd753: poly = 10'd326;
            10'd754: poly = 10'd652;
            10'd755: poly = 10'd273;
            10'd756: poly = 10'd546;
            10'd757: poly = 10'd77;
            10'd758: poly = 10'd154;
            10'd759: poly = 10'd308;
            10'd760: poly = 10'd616;
            10'd761: poly = 10'd217;
            10'd762: poly = 10'd434;
            10'd763: poly = 10'd868;
            10'd764: poly = 10'd705;
            10'd765: poly = 10'd395;
            10'd766: poly = 10'd790;
            10'd767: poly = 10'd549;
            10'd768: poly = 10'd67;
            10'd769: poly = 10'd134;
            10'd770: poly = 10'd268;
            10'd771: poly = 10'd536;
            10'd772: poly = 10'd57;
            10'd773: poly = 10'd114;
            10'd774: poly = 10'd228;
            10'd775: poly = 10'd456;
            10'd776: poly = 10'd912;
            10'd777: poly = 10'd809;
            10'd778: poly = 10'd603;
            10'd779: poly = 10'd191;
            10'd780: poly = 10'd382;
            10'd781: poly = 10'd764;
            10'd782: poly = 10'd497;
            10'd783: poly = 10'd994;
            10'd784: poly = 10'd973;
            10'd785: poly = 10'd915;
            10'd786: poly = 10'd815;
            10'd787: poly = 10'd599;
            10'd788: poly = 10'd167;
            10'd789: poly = 10'd334;
            10'd790: poly = 10'd668;
            10'd791: poly = 10'd305;
            10'd792: poly = 10'd610;
            10'd793: poly = 10'd205;
            10'd794: poly = 10'd410;
            10'd795: poly = 10'd820;
            10'd796: poly = 10'd609;
            10'd797: poly = 10'd203;
            10'd798: poly = 10'd406;
            10'd799: poly = 10'd812;
            10'd800: poly = 10'd593;
            10'd801: poly = 10'd171;
            10'd802: poly = 10'd342;
            10'd803: poly = 10'd684;
            10'd804: poly = 10'd337;
            10'd805: poly = 10'd674;
            10'd806: poly = 10'd333;
            10'd807: poly = 10'd666;
            10'd808: poly = 10'd317;
            10'd809: poly = 10'd634;
            10'd810: poly = 10'd253;
            10'd811: poly = 10'd506;
            10'd812: poly = 10'd1012;
            10'd813: poly = 10'd993;
            10'd814: poly = 10'd971;
            10'd815: poly = 10'd927;
            10'd816: poly = 10'd823;
            10'd817: poly = 10'd615;
            10'd818: poly = 10'd199;
            10'd819: poly = 10'd398;
            10'd820: poly = 10'd796;
            10'd821: poly = 10'd561;
            10'd822: poly = 10'd107;
            10'd823: poly = 10'd214;
            10'd824: poly = 10'd428;
            10'd825: poly = 10'd856;
            10'd826: poly = 10'd697;
            10'd827: poly = 10'd379;
            10'd828: poly = 10'd758;
            10'd829: poly = 10'd485;
            10'd830: poly = 10'd970;
            10'd831: poly = 10'd925;
            10'd832: poly = 10'd819;
            10'd833: poly = 10'd623;
            10'd834: poly = 10'd215;
            10'd835: poly = 10'd430;
            10'd836: poly = 10'd860;
            10'd837: poly = 10'd689;
            10'd838: poly = 10'd363;
            10'd839: poly = 10'd726;
            10'd840: poly = 10'd421;
            10'd841: poly = 10'd842;
            10'd842: poly = 10'd669;
            10'd843: poly = 10'd307;
            10'd844: poly = 10'd614;
            10'd845: poly = 10'd197;
            10'd846: poly = 10'd394;
            10'd847: poly = 10'd788;
            10'd848: poly = 10'd545;
            10'd849: poly = 10'd75;
            10'd850: poly = 10'd150;
            10'd851: poly = 10'd300;
            10'd852: poly = 10'd600;
            10'd853: poly = 10'd185;
            10'd854: poly = 10'd370;
            10'd855: poly = 10'd740;
            10'd856: poly = 10'd449;
            10'd857: poly = 10'd898;
            10'd858: poly = 10'd781;
            10'd859: poly = 10'd531;
            10'd860: poly = 10'd47;
            10'd861: poly = 10'd94;
            10'd862: poly = 10'd188;
            10'd863: poly = 10'd376;
            10'd864: poly = 10'd752;
            10'd865: poly = 10'd489;
            10'd866: poly = 10'd978;
            10'd867: poly = 10'd941;
            10'd868: poly = 10'd851;
            10'd869: poly = 10'd687;
            10'd870: poly = 10'd343;
            10'd871: poly = 10'd686;
            10'd872: poly = 10'd341;
            10'd873: poly = 10'd682;
            10'd874: poly = 10'd349;
            10'd875: poly = 10'd698;
            10'd876: poly = 10'd381;
            10'd877: poly = 10'd762;
            10'd878: poly = 10'd509;
            10'd879: poly = 10'd1018;
            10'd880: poly = 10'd1021;
            10'd881: poly = 10'd1011;
            10'd882: poly = 10'd1007;
            10'd883: poly = 10'd983;
            10'd884: poly = 10'd935;
            10'd885: poly = 10'd839;
            10'd886: poly = 10'd647;
            10'd887: poly = 10'd263;
            10'd888: poly = 10'd526;
            10'd889: poly = 10'd21;
            10'd890: poly = 10'd42;
            10'd891: poly = 10'd84;
            10'd892: poly = 10'd168;
            10'd893: poly = 10'd336;
            10'd894: poly = 10'd672;
            10'd895: poly = 10'd329;
            10'd896: poly = 10'd658;
            10'd897: poly = 10'd301;
            10'd898: poly = 10'd602;
            10'd899: poly = 10'd189;
            10'd900: poly = 10'd378;
            10'd901: poly = 10'd756;
            10'd902: poly = 10'd481;
            10'd903: poly = 10'd962;
            10'd904: poly = 10'd909;
            10'd905: poly = 10'd787;
            10'd906: poly = 10'd559;
            10'd907: poly = 10'd87;
            10'd908: poly = 10'd174;
            10'd909: poly = 10'd348;
            10'd910: poly = 10'd696;
            10'd911: poly = 10'd377;
            10'd912: poly = 10'd754;
            10'd913: poly = 10'd493;
            10'd914: poly = 10'd986;
            10'd915: poly = 10'd957;
            10'd916: poly = 10'd883;
            10'd917: poly = 10'd751;
            10'd918: poly = 10'd471;
            10'd919: poly = 10'd942;
            10'd920: poly = 10'd853;
            10'd921: poly = 10'd675;
            10'd922: poly = 10'd335;
            10'd923: poly = 10'd670;
            10'd924: poly = 10'd309;
            10'd925: poly = 10'd618;
            10'd926: poly = 10'd221;
            10'd927: poly = 10'd442;
            10'd928: poly = 10'd884;
            10'd929: poly = 10'd737;
            10'd930: poly = 10'd459;
            10'd931: poly = 10'd918;
            10'd932: poly = 10'd805;
            10'd933: poly = 10'd579;
            10'd934: poly = 10'd143;
            10'd935: poly = 10'd286;
            10'd936: poly = 10'd572;
            10'd937: poly = 10'd113;
            10'd938: poly = 10'd226;
            10'd939: poly = 10'd452;
            10'd940: poly = 10'd904;
            10'd941: poly = 10'd793;
            10'd942: poly = 10'd571;
            10'd943: poly = 10'd127;
            10'd944: poly = 10'd254;
            10'd945: poly = 10'd508;
            10'd946: poly = 10'd1016;
            10'd947: poly = 10'd1017;
            10'd948: poly = 10'd1019;
            10'd949: poly = 10'd1023;
            10'd950: poly = 10'd1015;
            10'd951: poly = 10'd999;
            10'd952: poly = 10'd967;
            10'd953: poly = 10'd903;
            10'd954: poly = 10'd775;
            10'd955: poly = 10'd519;
            10'd956: poly = 10'd7;
            10'd957: poly = 10'd14;
            10'd958: poly = 10'd28;
            10'd959: poly = 10'd56;
            10'd960: poly = 10'd112;
            10'd961: poly = 10'd224;
            10'd962: poly = 10'd448;
            10'd963: poly = 10'd896;
            10'd964: poly = 10'd777;
            10'd965: poly = 10'd539;
            10'd966: poly = 10'd63;
            10'd967: poly = 10'd126;
            10'd968: poly = 10'd252;
            10'd969: poly = 10'd504;
            10'd970: poly = 10'd1008;
            10'd971: poly = 10'd1001;
            10'd972: poly = 10'd987;
            10'd973: poly = 10'd959;
            10'd974: poly = 10'd887;
            10'd975: poly = 10'd743;
            10'd976: poly = 10'd455;
            10'd977: poly = 10'd910;
            10'd978: poly = 10'd789;
            10'd979: poly = 10'd547;
            10'd980: poly = 10'd79;
            10'd981: poly = 10'd158;
            10'd982: poly = 10'd316;
            10'd983: poly = 10'd632;
            10'd984: poly = 10'd249;
            10'd985: poly = 10'd498;
            10'd986: poly = 10'd996;
            10'd987: poly = 10'd961;
            10'd988: poly = 10'd907;
            10'd989: poly = 10'd799;
            10'd990: poly = 10'd567;
            10'd991: poly = 10'd103;
            10'd992: poly = 10'd206;
            10'd993: poly = 10'd412;
            10'd994: poly = 10'd824;
            10'd995: poly = 10'd633;
            10'd996: poly = 10'd251;
            10'd997: poly = 10'd502;
            10'd998: poly = 10'd1004;
            10'd999: poly = 10'd977;
            10'd1000: poly = 10'd939;
            10'd1001: poly = 10'd863;
            10'd1002: poly = 10'd695;
            10'd1003: poly = 10'd359;
            10'd1004: poly = 10'd718;
            10'd1005: poly = 10'd405;
            10'd1006: poly = 10'd810;
            10'd1007: poly = 10'd605;
            10'd1008: poly = 10'd179;
            10'd1009: poly = 10'd358;
            10'd1010: poly = 10'd716;
            10'd1011: poly = 10'd401;
            10'd1012: poly = 10'd802;
            10'd1013: poly = 10'd589;
            10'd1014: poly = 10'd147;
            10'd1015: poly = 10'd294;
            10'd1016: poly = 10'd588;
            10'd1017: poly = 10'd145;
            10'd1018: poly = 10'd290;
            10'd1019: poly = 10'd580;
            10'd1020: poly = 10'd129;
            10'd1021: poly = 10'd258;
            10'd1022: poly = 10'd516;
            default : poly = 10'd0;
        endcase
    end
endmodule

module GF_10_inv (
	input [9:0] poly,
	output reg [9:0] power
);
    always @* begin
        case(poly)
            10'd0: power = 10'd-1;
            10'd1: power = 10'd0;
            10'd2: power = 10'd1;
            10'd4: power = 10'd2;
            10'd8: power = 10'd3;
            10'd16: power = 10'd4;
            10'd32: power = 10'd5;
            10'd64: power = 10'd6;
            10'd128: power = 10'd7;
            10'd256: power = 10'd8;
            10'd512: power = 10'd9;
            10'd9: power = 10'd10;
            10'd18: power = 10'd11;
            10'd36: power = 10'd12;
            10'd72: power = 10'd13;
            10'd144: power = 10'd14;
            10'd288: power = 10'd15;
            10'd576: power = 10'd16;
            10'd137: power = 10'd17;
            10'd274: power = 10'd18;
            10'd548: power = 10'd19;
            10'd65: power = 10'd20;
            10'd130: power = 10'd21;
            10'd260: power = 10'd22;
            10'd520: power = 10'd23;
            10'd25: power = 10'd24;
            10'd50: power = 10'd25;
            10'd100: power = 10'd26;
            10'd200: power = 10'd27;
            10'd400: power = 10'd28;
            10'd800: power = 10'd29;
            10'd585: power = 10'd30;
            10'd155: power = 10'd31;
            10'd310: power = 10'd32;
            10'd620: power = 10'd33;
            10'd209: power = 10'd34;
            10'd418: power = 10'd35;
            10'd836: power = 10'd36;
            10'd641: power = 10'd37;
            10'd267: power = 10'd38;
            10'd534: power = 10'd39;
            10'd37: power = 10'd40;
            10'd74: power = 10'd41;
            10'd148: power = 10'd42;
            10'd296: power = 10'd43;
            10'd592: power = 10'd44;
            10'd169: power = 10'd45;
            10'd338: power = 10'd46;
            10'd676: power = 10'd47;
            10'd321: power = 10'd48;
            10'd642: power = 10'd49;
            10'd269: power = 10'd50;
            10'd538: power = 10'd51;
            10'd61: power = 10'd52;
            10'd122: power = 10'd53;
            10'd244: power = 10'd54;
            10'd488: power = 10'd55;
            10'd976: power = 10'd56;
            10'd937: power = 10'd57;
            10'd859: power = 10'd58;
            10'd703: power = 10'd59;
            10'd375: power = 10'd60;
            10'd750: power = 10'd61;
            10'd469: power = 10'd62;
            10'd938: power = 10'd63;
            10'd861: power = 10'd64;
            10'd691: power = 10'd65;
            10'd367: power = 10'd66;
            10'd734: power = 10'd67;
            10'd437: power = 10'd68;
            10'd874: power = 10'd69;
            10'd733: power = 10'd70;
            10'd435: power = 10'd71;
            10'd870: power = 10'd72;
            10'd709: power = 10'd73;
            10'd387: power = 10'd74;
            10'd774: power = 10'd75;
            10'd517: power = 10'd76;
            10'd3: power = 10'd77;
            10'd6: power = 10'd78;
            10'd12: power = 10'd79;
            10'd24: power = 10'd80;
            10'd48: power = 10'd81;
            10'd96: power = 10'd82;
            10'd192: power = 10'd83;
            10'd384: power = 10'd84;
            10'd768: power = 10'd85;
            10'd521: power = 10'd86;
            10'd27: power = 10'd87;
            10'd54: power = 10'd88;
            10'd108: power = 10'd89;
            10'd216: power = 10'd90;
            10'd432: power = 10'd91;
            10'd864: power = 10'd92;
            10'd713: power = 10'd93;
            10'd411: power = 10'd94;
            10'd822: power = 10'd95;
            10'd613: power = 10'd96;
            10'd195: power = 10'd97;
            10'd390: power = 10'd98;
            10'd780: power = 10'd99;
            10'd529: power = 10'd100;
            10'd43: power = 10'd101;
            10'd86: power = 10'd102;
            10'd172: power = 10'd103;
            10'd344: power = 10'd104;
            10'd688: power = 10'd105;
            10'd361: power = 10'd106;
            10'd722: power = 10'd107;
            10'd429: power = 10'd108;
            10'd858: power = 10'd109;
            10'd701: power = 10'd110;
            10'd371: power = 10'd111;
            10'd742: power = 10'd112;
            10'd453: power = 10'd113;
            10'd906: power = 10'd114;
            10'd797: power = 10'd115;
            10'd563: power = 10'd116;
            10'd111: power = 10'd117;
            10'd222: power = 10'd118;
            10'd444: power = 10'd119;
            10'd888: power = 10'd120;
            10'd761: power = 10'd121;
            10'd507: power = 10'd122;
            10'd1014: power = 10'd123;
            10'd997: power = 10'd124;
            10'd963: power = 10'd125;
            10'd911: power = 10'd126;
            10'd791: power = 10'd127;
            10'd551: power = 10'd128;
            10'd71: power = 10'd129;
            10'd142: power = 10'd130;
            10'd284: power = 10'd131;
            10'd568: power = 10'd132;
            10'd121: power = 10'd133;
            10'd242: power = 10'd134;
            10'd484: power = 10'd135;
            10'd968: power = 10'd136;
            10'd921: power = 10'd137;
            10'd827: power = 10'd138;
            10'd639: power = 10'd139;
            10'd247: power = 10'd140;
            10'd494: power = 10'd141;
            10'd988: power = 10'd142;
            10'd945: power = 10'd143;
            10'd875: power = 10'd144;
            10'd735: power = 10'd145;
            10'd439: power = 10'd146;
            10'd878: power = 10'd147;
            10'd725: power = 10'd148;
            10'd419: power = 10'd149;
            10'd838: power = 10'd150;
            10'd645: power = 10'd151;
            10'd259: power = 10'd152;
            10'd518: power = 10'd153;
            10'd5: power = 10'd154;
            10'd10: power = 10'd155;
            10'd20: power = 10'd156;
            10'd40: power = 10'd157;
            10'd80: power = 10'd158;
            10'd160: power = 10'd159;
            10'd320: power = 10'd160;
            10'd640: power = 10'd161;
            10'd265: power = 10'd162;
            10'd530: power = 10'd163;
            10'd45: power = 10'd164;
            10'd90: power = 10'd165;
            10'd180: power = 10'd166;
            10'd360: power = 10'd167;
            10'd720: power = 10'd168;
            10'd425: power = 10'd169;
            10'd850: power = 10'd170;
            10'd685: power = 10'd171;
            10'd339: power = 10'd172;
            10'd678: power = 10'd173;
            10'd325: power = 10'd174;
            10'd650: power = 10'd175;
            10'd285: power = 10'd176;
            10'd570: power = 10'd177;
            10'd125: power = 10'd178;
            10'd250: power = 10'd179;
            10'd500: power = 10'd180;
            10'd1000: power = 10'd181;
            10'd985: power = 10'd182;
            10'd955: power = 10'd183;
            10'd895: power = 10'd184;
            10'd759: power = 10'd185;
            10'd487: power = 10'd186;
            10'd974: power = 10'd187;
            10'd917: power = 10'd188;
            10'd803: power = 10'd189;
            10'd591: power = 10'd190;
            10'd151: power = 10'd191;
            10'd302: power = 10'd192;
            10'd604: power = 10'd193;
            10'd177: power = 10'd194;
            10'd354: power = 10'd195;
            10'd708: power = 10'd196;
            10'd385: power = 10'd197;
            10'd770: power = 10'd198;
            10'd525: power = 10'd199;
            10'd19: power = 10'd200;
            10'd38: power = 10'd201;
            10'd76: power = 10'd202;
            10'd152: power = 10'd203;
            10'd304: power = 10'd204;
            10'd608: power = 10'd205;
            10'd201: power = 10'd206;
            10'd402: power = 10'd207;
            10'd804: power = 10'd208;
            10'd577: power = 10'd209;
            10'd139: power = 10'd210;
            10'd278: power = 10'd211;
            10'd556: power = 10'd212;
            10'd81: power = 10'd213;
            10'd162: power = 10'd214;
            10'd324: power = 10'd215;
            10'd648: power = 10'd216;
            10'd281: power = 10'd217;
            10'd562: power = 10'd218;
            10'd109: power = 10'd219;
            10'd218: power = 10'd220;
            10'd436: power = 10'd221;
            10'd872: power = 10'd222;
            10'd729: power = 10'd223;
            10'd443: power = 10'd224;
            10'd886: power = 10'd225;
            10'd741: power = 10'd226;
            10'd451: power = 10'd227;
            10'd902: power = 10'd228;
            10'd773: power = 10'd229;
            10'd515: power = 10'd230;
            10'd15: power = 10'd231;
            10'd30: power = 10'd232;
            10'd60: power = 10'd233;
            10'd120: power = 10'd234;
            10'd240: power = 10'd235;
            10'd480: power = 10'd236;
            10'd960: power = 10'd237;
            10'd905: power = 10'd238;
            10'd795: power = 10'd239;
            10'd575: power = 10'd240;
            10'd119: power = 10'd241;
            10'd238: power = 10'd242;
            10'd476: power = 10'd243;
            10'd952: power = 10'd244;
            10'd889: power = 10'd245;
            10'd763: power = 10'd246;
            10'd511: power = 10'd247;
            10'd1022: power = 10'd248;
            10'd1013: power = 10'd249;
            10'd995: power = 10'd250;
            10'd975: power = 10'd251;
            10'd919: power = 10'd252;
            10'd807: power = 10'd253;
            10'd583: power = 10'd254;
            10'd135: power = 10'd255;
            10'd270: power = 10'd256;
            10'd540: power = 10'd257;
            10'd49: power = 10'd258;
            10'd98: power = 10'd259;
            10'd196: power = 10'd260;
            10'd392: power = 10'd261;
            10'd784: power = 10'd262;
            10'd553: power = 10'd263;
            10'd91: power = 10'd264;
            10'd182: power = 10'd265;
            10'd364: power = 10'd266;
            10'd728: power = 10'd267;
            10'd441: power = 10'd268;
            10'd882: power = 10'd269;
            10'd749: power = 10'd270;
            10'd467: power = 10'd271;
            10'd934: power = 10'd272;
            10'd837: power = 10'd273;
            10'd643: power = 10'd274;
            10'd271: power = 10'd275;
            10'd542: power = 10'd276;
            10'd53: power = 10'd277;
            10'd106: power = 10'd278;
            10'd212: power = 10'd279;
            10'd424: power = 10'd280;
            10'd848: power = 10'd281;
            10'd681: power = 10'd282;
            10'd347: power = 10'd283;
            10'd694: power = 10'd284;
            10'd357: power = 10'd285;
            10'd714: power = 10'd286;
            10'd413: power = 10'd287;
            10'd826: power = 10'd288;
            10'd637: power = 10'd289;
            10'd243: power = 10'd290;
            10'd486: power = 10'd291;
            10'd972: power = 10'd292;
            10'd913: power = 10'd293;
            10'd811: power = 10'd294;
            10'd607: power = 10'd295;
            10'd183: power = 10'd296;
            10'd366: power = 10'd297;
            10'd732: power = 10'd298;
            10'd433: power = 10'd299;
            10'd866: power = 10'd300;
            10'd717: power = 10'd301;
            10'd403: power = 10'd302;
            10'd806: power = 10'd303;
            10'd581: power = 10'd304;
            10'd131: power = 10'd305;
            10'd262: power = 10'd306;
            10'd524: power = 10'd307;
            10'd17: power = 10'd308;
            10'd34: power = 10'd309;
            10'd68: power = 10'd310;
            10'd136: power = 10'd311;
            10'd272: power = 10'd312;
            10'd544: power = 10'd313;
            10'd73: power = 10'd314;
            10'd146: power = 10'd315;
            10'd292: power = 10'd316;
            10'd584: power = 10'd317;
            10'd153: power = 10'd318;
            10'd306: power = 10'd319;
            10'd612: power = 10'd320;
            10'd193: power = 10'd321;
            10'd386: power = 10'd322;
            10'd772: power = 10'd323;
            10'd513: power = 10'd324;
            10'd11: power = 10'd325;
            10'd22: power = 10'd326;
            10'd44: power = 10'd327;
            10'd88: power = 10'd328;
            10'd176: power = 10'd329;
            10'd352: power = 10'd330;
            10'd704: power = 10'd331;
            10'd393: power = 10'd332;
            10'd786: power = 10'd333;
            10'd557: power = 10'd334;
            10'd83: power = 10'd335;
            10'd166: power = 10'd336;
            10'd332: power = 10'd337;
            10'd664: power = 10'd338;
            10'd313: power = 10'd339;
            10'd626: power = 10'd340;
            10'd237: power = 10'd341;
            10'd474: power = 10'd342;
            10'd948: power = 10'd343;
            10'd865: power = 10'd344;
            10'd715: power = 10'd345;
            10'd415: power = 10'd346;
            10'd830: power = 10'd347;
            10'd629: power = 10'd348;
            10'd227: power = 10'd349;
            10'd454: power = 10'd350;
            10'd908: power = 10'd351;
            10'd785: power = 10'd352;
            10'd555: power = 10'd353;
            10'd95: power = 10'd354;
            10'd190: power = 10'd355;
            10'd380: power = 10'd356;
            10'd760: power = 10'd357;
            10'd505: power = 10'd358;
            10'd1010: power = 10'd359;
            10'd1005: power = 10'd360;
            10'd979: power = 10'd361;
            10'd943: power = 10'd362;
            10'd855: power = 10'd363;
            10'd679: power = 10'd364;
            10'd327: power = 10'd365;
            10'd654: power = 10'd366;
            10'd277: power = 10'd367;
            10'd554: power = 10'd368;
            10'd93: power = 10'd369;
            10'd186: power = 10'd370;
            10'd372: power = 10'd371;
            10'd744: power = 10'd372;
            10'd473: power = 10'd373;
            10'd946: power = 10'd374;
            10'd877: power = 10'd375;
            10'd723: power = 10'd376;
            10'd431: power = 10'd377;
            10'd862: power = 10'd378;
            10'd693: power = 10'd379;
            10'd355: power = 10'd380;
            10'd710: power = 10'd381;
            10'd389: power = 10'd382;
            10'd778: power = 10'd383;
            10'd541: power = 10'd384;
            10'd51: power = 10'd385;
            10'd102: power = 10'd386;
            10'd204: power = 10'd387;
            10'd408: power = 10'd388;
            10'd816: power = 10'd389;
            10'd617: power = 10'd390;
            10'd219: power = 10'd391;
            10'd438: power = 10'd392;
            10'd876: power = 10'd393;
            10'd721: power = 10'd394;
            10'd427: power = 10'd395;
            10'd854: power = 10'd396;
            10'd677: power = 10'd397;
            10'd323: power = 10'd398;
            10'd646: power = 10'd399;
            10'd261: power = 10'd400;
            10'd522: power = 10'd401;
            10'd29: power = 10'd402;
            10'd58: power = 10'd403;
            10'd116: power = 10'd404;
            10'd232: power = 10'd405;
            10'd464: power = 10'd406;
            10'd928: power = 10'd407;
            10'd841: power = 10'd408;
            10'd667: power = 10'd409;
            10'd319: power = 10'd410;
            10'd638: power = 10'd411;
            10'd245: power = 10'd412;
            10'd490: power = 10'd413;
            10'd980: power = 10'd414;
            10'd929: power = 10'd415;
            10'd843: power = 10'd416;
            10'd671: power = 10'd417;
            10'd311: power = 10'd418;
            10'd622: power = 10'd419;
            10'd213: power = 10'd420;
            10'd426: power = 10'd421;
            10'd852: power = 10'd422;
            10'd673: power = 10'd423;
            10'd331: power = 10'd424;
            10'd662: power = 10'd425;
            10'd293: power = 10'd426;
            10'd586: power = 10'd427;
            10'd157: power = 10'd428;
            10'd314: power = 10'd429;
            10'd628: power = 10'd430;
            10'd225: power = 10'd431;
            10'd450: power = 10'd432;
            10'd900: power = 10'd433;
            10'd769: power = 10'd434;
            10'd523: power = 10'd435;
            10'd31: power = 10'd436;
            10'd62: power = 10'd437;
            10'd124: power = 10'd438;
            10'd248: power = 10'd439;
            10'd496: power = 10'd440;
            10'd992: power = 10'd441;
            10'd969: power = 10'd442;
            10'd923: power = 10'd443;
            10'd831: power = 10'd444;
            10'd631: power = 10'd445;
            10'd231: power = 10'd446;
            10'd462: power = 10'd447;
            10'd924: power = 10'd448;
            10'd817: power = 10'd449;
            10'd619: power = 10'd450;
            10'd223: power = 10'd451;
            10'd446: power = 10'd452;
            10'd892: power = 10'd453;
            10'd753: power = 10'd454;
            10'd491: power = 10'd455;
            10'd982: power = 10'd456;
            10'd933: power = 10'd457;
            10'd835: power = 10'd458;
            10'd655: power = 10'd459;
            10'd279: power = 10'd460;
            10'd558: power = 10'd461;
            10'd85: power = 10'd462;
            10'd170: power = 10'd463;
            10'd340: power = 10'd464;
            10'd680: power = 10'd465;
            10'd345: power = 10'd466;
            10'd690: power = 10'd467;
            10'd365: power = 10'd468;
            10'd730: power = 10'd469;
            10'd445: power = 10'd470;
            10'd890: power = 10'd471;
            10'd765: power = 10'd472;
            10'd499: power = 10'd473;
            10'd998: power = 10'd474;
            10'd965: power = 10'd475;
            10'd899: power = 10'd476;
            10'd783: power = 10'd477;
            10'd535: power = 10'd478;
            10'd39: power = 10'd479;
            10'd78: power = 10'd480;
            10'd156: power = 10'd481;
            10'd312: power = 10'd482;
            10'd624: power = 10'd483;
            10'd233: power = 10'd484;
            10'd466: power = 10'd485;
            10'd932: power = 10'd486;
            10'd833: power = 10'd487;
            10'd651: power = 10'd488;
            10'd287: power = 10'd489;
            10'd574: power = 10'd490;
            10'd117: power = 10'd491;
            10'd234: power = 10'd492;
            10'd468: power = 10'd493;
            10'd936: power = 10'd494;
            10'd857: power = 10'd495;
            10'd699: power = 10'd496;
            10'd383: power = 10'd497;
            10'd766: power = 10'd498;
            10'd501: power = 10'd499;
            10'd1002: power = 10'd500;
            10'd989: power = 10'd501;
            10'd947: power = 10'd502;
            10'd879: power = 10'd503;
            10'd727: power = 10'd504;
            10'd423: power = 10'd505;
            10'd846: power = 10'd506;
            10'd661: power = 10'd507;
            10'd291: power = 10'd508;
            10'd582: power = 10'd509;
            10'd133: power = 10'd510;
            10'd266: power = 10'd511;
            10'd532: power = 10'd512;
            10'd33: power = 10'd513;
            10'd66: power = 10'd514;
            10'd132: power = 10'd515;
            10'd264: power = 10'd516;
            10'd528: power = 10'd517;
            10'd41: power = 10'd518;
            10'd82: power = 10'd519;
            10'd164: power = 10'd520;
            10'd328: power = 10'd521;
            10'd656: power = 10'd522;
            10'd297: power = 10'd523;
            10'd594: power = 10'd524;
            10'd173: power = 10'd525;
            10'd346: power = 10'd526;
            10'd692: power = 10'd527;
            10'd353: power = 10'd528;
            10'd706: power = 10'd529;
            10'd397: power = 10'd530;
            10'd794: power = 10'd531;
            10'd573: power = 10'd532;
            10'd115: power = 10'd533;
            10'd230: power = 10'd534;
            10'd460: power = 10'd535;
            10'd920: power = 10'd536;
            10'd825: power = 10'd537;
            10'd635: power = 10'd538;
            10'd255: power = 10'd539;
            10'd510: power = 10'd540;
            10'd1020: power = 10'd541;
            10'd1009: power = 10'd542;
            10'd1003: power = 10'd543;
            10'd991: power = 10'd544;
            10'd951: power = 10'd545;
            10'd871: power = 10'd546;
            10'd711: power = 10'd547;
            10'd391: power = 10'd548;
            10'd782: power = 10'd549;
            10'd533: power = 10'd550;
            10'd35: power = 10'd551;
            10'd70: power = 10'd552;
            10'd140: power = 10'd553;
            10'd280: power = 10'd554;
            10'd560: power = 10'd555;
            10'd105: power = 10'd556;
            10'd210: power = 10'd557;
            10'd420: power = 10'd558;
            10'd840: power = 10'd559;
            10'd665: power = 10'd560;
            10'd315: power = 10'd561;
            10'd630: power = 10'd562;
            10'd229: power = 10'd563;
            10'd458: power = 10'd564;
            10'd916: power = 10'd565;
            10'd801: power = 10'd566;
            10'd587: power = 10'd567;
            10'd159: power = 10'd568;
            10'd318: power = 10'd569;
            10'd636: power = 10'd570;
            10'd241: power = 10'd571;
            10'd482: power = 10'd572;
            10'd964: power = 10'd573;
            10'd897: power = 10'd574;
            10'd779: power = 10'd575;
            10'd543: power = 10'd576;
            10'd55: power = 10'd577;
            10'd110: power = 10'd578;
            10'd220: power = 10'd579;
            10'd440: power = 10'd580;
            10'd880: power = 10'd581;
            10'd745: power = 10'd582;
            10'd475: power = 10'd583;
            10'd950: power = 10'd584;
            10'd869: power = 10'd585;
            10'd707: power = 10'd586;
            10'd399: power = 10'd587;
            10'd798: power = 10'd588;
            10'd565: power = 10'd589;
            10'd99: power = 10'd590;
            10'd198: power = 10'd591;
            10'd396: power = 10'd592;
            10'd792: power = 10'd593;
            10'd569: power = 10'd594;
            10'd123: power = 10'd595;
            10'd246: power = 10'd596;
            10'd492: power = 10'd597;
            10'd984: power = 10'd598;
            10'd953: power = 10'd599;
            10'd891: power = 10'd600;
            10'd767: power = 10'd601;
            10'd503: power = 10'd602;
            10'd1006: power = 10'd603;
            10'd981: power = 10'd604;
            10'd931: power = 10'd605;
            10'd847: power = 10'd606;
            10'd663: power = 10'd607;
            10'd295: power = 10'd608;
            10'd590: power = 10'd609;
            10'd149: power = 10'd610;
            10'd298: power = 10'd611;
            10'd596: power = 10'd612;
            10'd161: power = 10'd613;
            10'd322: power = 10'd614;
            10'd644: power = 10'd615;
            10'd257: power = 10'd616;
            10'd514: power = 10'd617;
            10'd13: power = 10'd618;
            10'd26: power = 10'd619;
            10'd52: power = 10'd620;
            10'd104: power = 10'd621;
            10'd208: power = 10'd622;
            10'd416: power = 10'd623;
            10'd832: power = 10'd624;
            10'd649: power = 10'd625;
            10'd283: power = 10'd626;
            10'd566: power = 10'd627;
            10'd101: power = 10'd628;
            10'd202: power = 10'd629;
            10'd404: power = 10'd630;
            10'd808: power = 10'd631;
            10'd601: power = 10'd632;
            10'd187: power = 10'd633;
            10'd374: power = 10'd634;
            10'd748: power = 10'd635;
            10'd465: power = 10'd636;
            10'd930: power = 10'd637;
            10'd845: power = 10'd638;
            10'd659: power = 10'd639;
            10'd303: power = 10'd640;
            10'd606: power = 10'd641;
            10'd181: power = 10'd642;
            10'd362: power = 10'd643;
            10'd724: power = 10'd644;
            10'd417: power = 10'd645;
            10'd834: power = 10'd646;
            10'd653: power = 10'd647;
            10'd275: power = 10'd648;
            10'd550: power = 10'd649;
            10'd69: power = 10'd650;
            10'd138: power = 10'd651;
            10'd276: power = 10'd652;
            10'd552: power = 10'd653;
            10'd89: power = 10'd654;
            10'd178: power = 10'd655;
            10'd356: power = 10'd656;
            10'd712: power = 10'd657;
            10'd409: power = 10'd658;
            10'd818: power = 10'd659;
            10'd621: power = 10'd660;
            10'd211: power = 10'd661;
            10'd422: power = 10'd662;
            10'd844: power = 10'd663;
            10'd657: power = 10'd664;
            10'd299: power = 10'd665;
            10'd598: power = 10'd666;
            10'd165: power = 10'd667;
            10'd330: power = 10'd668;
            10'd660: power = 10'd669;
            10'd289: power = 10'd670;
            10'd578: power = 10'd671;
            10'd141: power = 10'd672;
            10'd282: power = 10'd673;
            10'd564: power = 10'd674;
            10'd97: power = 10'd675;
            10'd194: power = 10'd676;
            10'd388: power = 10'd677;
            10'd776: power = 10'd678;
            10'd537: power = 10'd679;
            10'd59: power = 10'd680;
            10'd118: power = 10'd681;
            10'd236: power = 10'd682;
            10'd472: power = 10'd683;
            10'd944: power = 10'd684;
            10'd873: power = 10'd685;
            10'd731: power = 10'd686;
            10'd447: power = 10'd687;
            10'd894: power = 10'd688;
            10'd757: power = 10'd689;
            10'd483: power = 10'd690;
            10'd966: power = 10'd691;
            10'd901: power = 10'd692;
            10'd771: power = 10'd693;
            10'd527: power = 10'd694;
            10'd23: power = 10'd695;
            10'd46: power = 10'd696;
            10'd92: power = 10'd697;
            10'd184: power = 10'd698;
            10'd368: power = 10'd699;
            10'd736: power = 10'd700;
            10'd457: power = 10'd701;
            10'd914: power = 10'd702;
            10'd813: power = 10'd703;
            10'd595: power = 10'd704;
            10'd175: power = 10'd705;
            10'd350: power = 10'd706;
            10'd700: power = 10'd707;
            10'd369: power = 10'd708;
            10'd738: power = 10'd709;
            10'd461: power = 10'd710;
            10'd922: power = 10'd711;
            10'd829: power = 10'd712;
            10'd627: power = 10'd713;
            10'd239: power = 10'd714;
            10'd478: power = 10'd715;
            10'd956: power = 10'd716;
            10'd881: power = 10'd717;
            10'd747: power = 10'd718;
            10'd479: power = 10'd719;
            10'd958: power = 10'd720;
            10'd885: power = 10'd721;
            10'd739: power = 10'd722;
            10'd463: power = 10'd723;
            10'd926: power = 10'd724;
            10'd821: power = 10'd725;
            10'd611: power = 10'd726;
            10'd207: power = 10'd727;
            10'd414: power = 10'd728;
            10'd828: power = 10'd729;
            10'd625: power = 10'd730;
            10'd235: power = 10'd731;
            10'd470: power = 10'd732;
            10'd940: power = 10'd733;
            10'd849: power = 10'd734;
            10'd683: power = 10'd735;
            10'd351: power = 10'd736;
            10'd702: power = 10'd737;
            10'd373: power = 10'd738;
            10'd746: power = 10'd739;
            10'd477: power = 10'd740;
            10'd954: power = 10'd741;
            10'd893: power = 10'd742;
            10'd755: power = 10'd743;
            10'd495: power = 10'd744;
            10'd990: power = 10'd745;
            10'd949: power = 10'd746;
            10'd867: power = 10'd747;
            10'd719: power = 10'd748;
            10'd407: power = 10'd749;
            10'd814: power = 10'd750;
            10'd597: power = 10'd751;
            10'd163: power = 10'd752;
            10'd326: power = 10'd753;
            10'd652: power = 10'd754;
            10'd273: power = 10'd755;
            10'd546: power = 10'd756;
            10'd77: power = 10'd757;
            10'd154: power = 10'd758;
            10'd308: power = 10'd759;
            10'd616: power = 10'd760;
            10'd217: power = 10'd761;
            10'd434: power = 10'd762;
            10'd868: power = 10'd763;
            10'd705: power = 10'd764;
            10'd395: power = 10'd765;
            10'd790: power = 10'd766;
            10'd549: power = 10'd767;
            10'd67: power = 10'd768;
            10'd134: power = 10'd769;
            10'd268: power = 10'd770;
            10'd536: power = 10'd771;
            10'd57: power = 10'd772;
            10'd114: power = 10'd773;
            10'd228: power = 10'd774;
            10'd456: power = 10'd775;
            10'd912: power = 10'd776;
            10'd809: power = 10'd777;
            10'd603: power = 10'd778;
            10'd191: power = 10'd779;
            10'd382: power = 10'd780;
            10'd764: power = 10'd781;
            10'd497: power = 10'd782;
            10'd994: power = 10'd783;
            10'd973: power = 10'd784;
            10'd915: power = 10'd785;
            10'd815: power = 10'd786;
            10'd599: power = 10'd787;
            10'd167: power = 10'd788;
            10'd334: power = 10'd789;
            10'd668: power = 10'd790;
            10'd305: power = 10'd791;
            10'd610: power = 10'd792;
            10'd205: power = 10'd793;
            10'd410: power = 10'd794;
            10'd820: power = 10'd795;
            10'd609: power = 10'd796;
            10'd203: power = 10'd797;
            10'd406: power = 10'd798;
            10'd812: power = 10'd799;
            10'd593: power = 10'd800;
            10'd171: power = 10'd801;
            10'd342: power = 10'd802;
            10'd684: power = 10'd803;
            10'd337: power = 10'd804;
            10'd674: power = 10'd805;
            10'd333: power = 10'd806;
            10'd666: power = 10'd807;
            10'd317: power = 10'd808;
            10'd634: power = 10'd809;
            10'd253: power = 10'd810;
            10'd506: power = 10'd811;
            10'd1012: power = 10'd812;
            10'd993: power = 10'd813;
            10'd971: power = 10'd814;
            10'd927: power = 10'd815;
            10'd823: power = 10'd816;
            10'd615: power = 10'd817;
            10'd199: power = 10'd818;
            10'd398: power = 10'd819;
            10'd796: power = 10'd820;
            10'd561: power = 10'd821;
            10'd107: power = 10'd822;
            10'd214: power = 10'd823;
            10'd428: power = 10'd824;
            10'd856: power = 10'd825;
            10'd697: power = 10'd826;
            10'd379: power = 10'd827;
            10'd758: power = 10'd828;
            10'd485: power = 10'd829;
            10'd970: power = 10'd830;
            10'd925: power = 10'd831;
            10'd819: power = 10'd832;
            10'd623: power = 10'd833;
            10'd215: power = 10'd834;
            10'd430: power = 10'd835;
            10'd860: power = 10'd836;
            10'd689: power = 10'd837;
            10'd363: power = 10'd838;
            10'd726: power = 10'd839;
            10'd421: power = 10'd840;
            10'd842: power = 10'd841;
            10'd669: power = 10'd842;
            10'd307: power = 10'd843;
            10'd614: power = 10'd844;
            10'd197: power = 10'd845;
            10'd394: power = 10'd846;
            10'd788: power = 10'd847;
            10'd545: power = 10'd848;
            10'd75: power = 10'd849;
            10'd150: power = 10'd850;
            10'd300: power = 10'd851;
            10'd600: power = 10'd852;
            10'd185: power = 10'd853;
            10'd370: power = 10'd854;
            10'd740: power = 10'd855;
            10'd449: power = 10'd856;
            10'd898: power = 10'd857;
            10'd781: power = 10'd858;
            10'd531: power = 10'd859;
            10'd47: power = 10'd860;
            10'd94: power = 10'd861;
            10'd188: power = 10'd862;
            10'd376: power = 10'd863;
            10'd752: power = 10'd864;
            10'd489: power = 10'd865;
            10'd978: power = 10'd866;
            10'd941: power = 10'd867;
            10'd851: power = 10'd868;
            10'd687: power = 10'd869;
            10'd343: power = 10'd870;
            10'd686: power = 10'd871;
            10'd341: power = 10'd872;
            10'd682: power = 10'd873;
            10'd349: power = 10'd874;
            10'd698: power = 10'd875;
            10'd381: power = 10'd876;
            10'd762: power = 10'd877;
            10'd509: power = 10'd878;
            10'd1018: power = 10'd879;
            10'd1021: power = 10'd880;
            10'd1011: power = 10'd881;
            10'd1007: power = 10'd882;
            10'd983: power = 10'd883;
            10'd935: power = 10'd884;
            10'd839: power = 10'd885;
            10'd647: power = 10'd886;
            10'd263: power = 10'd887;
            10'd526: power = 10'd888;
            10'd21: power = 10'd889;
            10'd42: power = 10'd890;
            10'd84: power = 10'd891;
            10'd168: power = 10'd892;
            10'd336: power = 10'd893;
            10'd672: power = 10'd894;
            10'd329: power = 10'd895;
            10'd658: power = 10'd896;
            10'd301: power = 10'd897;
            10'd602: power = 10'd898;
            10'd189: power = 10'd899;
            10'd378: power = 10'd900;
            10'd756: power = 10'd901;
            10'd481: power = 10'd902;
            10'd962: power = 10'd903;
            10'd909: power = 10'd904;
            10'd787: power = 10'd905;
            10'd559: power = 10'd906;
            10'd87: power = 10'd907;
            10'd174: power = 10'd908;
            10'd348: power = 10'd909;
            10'd696: power = 10'd910;
            10'd377: power = 10'd911;
            10'd754: power = 10'd912;
            10'd493: power = 10'd913;
            10'd986: power = 10'd914;
            10'd957: power = 10'd915;
            10'd883: power = 10'd916;
            10'd751: power = 10'd917;
            10'd471: power = 10'd918;
            10'd942: power = 10'd919;
            10'd853: power = 10'd920;
            10'd675: power = 10'd921;
            10'd335: power = 10'd922;
            10'd670: power = 10'd923;
            10'd309: power = 10'd924;
            10'd618: power = 10'd925;
            10'd221: power = 10'd926;
            10'd442: power = 10'd927;
            10'd884: power = 10'd928;
            10'd737: power = 10'd929;
            10'd459: power = 10'd930;
            10'd918: power = 10'd931;
            10'd805: power = 10'd932;
            10'd579: power = 10'd933;
            10'd143: power = 10'd934;
            10'd286: power = 10'd935;
            10'd572: power = 10'd936;
            10'd113: power = 10'd937;
            10'd226: power = 10'd938;
            10'd452: power = 10'd939;
            10'd904: power = 10'd940;
            10'd793: power = 10'd941;
            10'd571: power = 10'd942;
            10'd127: power = 10'd943;
            10'd254: power = 10'd944;
            10'd508: power = 10'd945;
            10'd1016: power = 10'd946;
            10'd1017: power = 10'd947;
            10'd1019: power = 10'd948;
            10'd1023: power = 10'd949;
            10'd1015: power = 10'd950;
            10'd999: power = 10'd951;
            10'd967: power = 10'd952;
            10'd903: power = 10'd953;
            10'd775: power = 10'd954;
            10'd519: power = 10'd955;
            10'd7: power = 10'd956;
            10'd14: power = 10'd957;
            10'd28: power = 10'd958;
            10'd56: power = 10'd959;
            10'd112: power = 10'd960;
            10'd224: power = 10'd961;
            10'd448: power = 10'd962;
            10'd896: power = 10'd963;
            10'd777: power = 10'd964;
            10'd539: power = 10'd965;
            10'd63: power = 10'd966;
            10'd126: power = 10'd967;
            10'd252: power = 10'd968;
            10'd504: power = 10'd969;
            10'd1008: power = 10'd970;
            10'd1001: power = 10'd971;
            10'd987: power = 10'd972;
            10'd959: power = 10'd973;
            10'd887: power = 10'd974;
            10'd743: power = 10'd975;
            10'd455: power = 10'd976;
            10'd910: power = 10'd977;
            10'd789: power = 10'd978;
            10'd547: power = 10'd979;
            10'd79: power = 10'd980;
            10'd158: power = 10'd981;
            10'd316: power = 10'd982;
            10'd632: power = 10'd983;
            10'd249: power = 10'd984;
            10'd498: power = 10'd985;
            10'd996: power = 10'd986;
            10'd961: power = 10'd987;
            10'd907: power = 10'd988;
            10'd799: power = 10'd989;
            10'd567: power = 10'd990;
            10'd103: power = 10'd991;
            10'd206: power = 10'd992;
            10'd412: power = 10'd993;
            10'd824: power = 10'd994;
            10'd633: power = 10'd995;
            10'd251: power = 10'd996;
            10'd502: power = 10'd997;
            10'd1004: power = 10'd998;
            10'd977: power = 10'd999;
            10'd939: power = 10'd1000;
            10'd863: power = 10'd1001;
            10'd695: power = 10'd1002;
            10'd359: power = 10'd1003;
            10'd718: power = 10'd1004;
            10'd405: power = 10'd1005;
            10'd810: power = 10'd1006;
            10'd605: power = 10'd1007;
            10'd179: power = 10'd1008;
            10'd358: power = 10'd1009;
            10'd716: power = 10'd1010;
            10'd401: power = 10'd1011;
            10'd802: power = 10'd1012;
            10'd589: power = 10'd1013;
            10'd147: power = 10'd1014;
            10'd294: power = 10'd1015;
            10'd588: power = 10'd1016;
            10'd145: power = 10'd1017;
            10'd290: power = 10'd1018;
            10'd580: power = 10'd1019;
            10'd129: power = 10'd1020;
            10'd258: power = 10'd1021;
            10'd516: power = 10'd1022;
            default: power = 10'd1023;
        endcase
    end
endmodule